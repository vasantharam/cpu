`include "eth_defs.vh"
module eth_rx_driver(rx_drv_rd_data, rx_drv_rd_valid, rx_drv_rd_ready, clk, rst);

endmodule
