`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    17:53:34 10/24/2020 
// Design Name: 
// Module Name:    noc_defs 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////


`define ST_NOC_IDLE 0
`define ST_NOC_WR_PORT0_RESPOND 1
`define ST_NOC_WR_PORT1_RESPOND 2
`define ST_NOC_RD_PORT0_RESPOND 3
`define ST_NOC_RD_PORT1_RESPOND 4
`define ST_NOC_RD_PORT2_RESPOND 5
